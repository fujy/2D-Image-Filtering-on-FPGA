----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:53:52 11/05/2015 
-- Design Name: 
-- Module Name:    FlipFlop - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FlipFlop is

generic (Bus_Width : integer := 8);
    Port (D: IN STD_LOGIC_VECTOR (Bus_Width-1 downto 0);
			 Q: OUT STD_LOGIC_VECTOR (Bus_Width-1 downto 0);
			 CLK: IN STD_LOGIC;
			 EN: IN STD_LOGIC;
			 RESET: IN STD_LOGIC);
end FlipFlop;

architecture Behavioral of FlipFlop is

signal temp : STD_LOGIC_VECTOR (Bus_Width-1 downto 0) := (others => '0');

begin

MsCV_demo: process (clk,reset)
begin

	if (reset ='1') then temp <= (others => '0');
	elsif rising_edge(clk)
	then
		if ( en = '1') then
			temp <= D;
		else
			temp <= (others => '0');
		end if;
	end if;

end process MsCV_demo;

Q <= temp;

end Behavioral;

